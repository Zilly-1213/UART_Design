`define VLD_DATA_WIDTH 8